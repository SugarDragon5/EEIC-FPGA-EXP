`include "module/xorshift.v"
`include "module/distance.v"
`include "module/seg7.sv"
`include "module/swap.sv"
`include "module/swap_adjacent.sv"
`include "module/graph.sv"
`include "module/tsp.sv"
`include "module/TSPTop_wrap.sv"
