`include "xorshift.v"
`include "distance.v"
`include "seg7.sv"
`include "swap.sv"
`include "graph.sv"
`include "tsp.sv"
`include "TSPTop_wrap.sv"